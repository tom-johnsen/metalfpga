// EXPECT=PASS
// Test: Concatenation edge cases
// Feature: Empty concat, single element, nested replication
// Expected: May fail - edge case concatenation

module test_concatenation_edge;
  reg [7:0] a, b, c;
  wire [7:0] single;
  wire [31:0] nested_rep;
  wire [15:0] mixed;

  assign single = {a};  // Single element concat
  assign nested_rep = {4{{2{a}}}};  // Nested replication: 4 copies of (2 copies of a)
  assign mixed = {2{a, b[3:0]}};  // Replicate concatenation

  initial begin
    a = 8'hAA;
    b = 8'h55;
  end
endmodule
