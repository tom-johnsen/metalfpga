// EXPECT=PASS
// Test: supply1 net type (constant 1)
// Feature: Power/ground nets
// Expected: Should fail - supply nets not yet implemented

module test_net_supply1(
  output supply1 vdd
);
  // supply1 is always driven to logic 1 with supply strength
endmodule
