// EXPECT=PASS
// Test: Gate array instantiation
// Feature: Gate-level primitives
// Expected: Should fail - gate primitives not yet implemented

module test_gate_array(input [3:0] a, input [3:0] b, output [3:0] y);
  and g[3:0](y, a, b);  // 4 parallel AND gates
endmodule
