// EXPECT=PASS
module comb_loop;
  wire a;
  wire b;

  assign a = b;
  assign b = a;
endmodule
