module negedge_ff(input clk, d, output reg q);
  always @(negedge clk) q <= d;
endmodule
