// EXPECT=PASS
// Test: Array of tristate buffers
// Feature: Gate arrays with tristate
// Expected: Should fail - tristate gate arrays not yet implemented

module test_tristate_array(
  input [7:0] data,
  input [7:0] enable,
  output [7:0] bus
);
  bufif1 buf_array[7:0](bus, data, enable);
  // 8 parallel tristate buffers, each controlled independently
endmodule
