// EXPECT=PASS
// Test: wand net type (wired-AND)
// Feature: Net types with implicit logic
// Expected: Should fail - wand not yet implemented

module test_net_wand(
  input a,
  input b,
  output wand y  // Wired-AND: y = a & b when both drive
);
  assign y = a;
  assign y = b;  // Multiple drivers on wand net
endmodule
