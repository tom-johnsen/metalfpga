// EXPECT=PASS
// Test: triand net type
// Feature: Tristate with wired-AND resolution
// Expected: Should fail - triand not yet implemented

module test_net_triand(
  input [7:0] data_a,
  input [7:0] data_b,
  input enable_a,
  input enable_b,
  output triand [7:0] bus
);
  assign bus = enable_a ? data_a : 8'bz;
  assign bus = enable_b ? data_b : 8'bz;
  // When both enabled, result is data_a & data_b
  // When one enabled, result is that data
  // When neither enabled, result is z
endmodule
