// EXPECT=PASS
// Test: $fopen, $fclose file operations
// Feature: File handle operations

module test_system_fopen;
  integer fd;

  initial begin
    fd = $fopen("output.txt", "w");   // Open for write
    if (fd)
      $fclose(fd);

    fd = $fopen("input.txt", "r");    // Open for read
    if (fd)
      $fclose(fd);

    fd = $fopen("append.txt", "a");   // Open for append
    if (fd)
      $fclose(fd);
  end
endmodule
