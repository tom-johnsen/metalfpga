// Shared definitions for include tests.
